package testb_pkg;
import uvm_pkg::*;
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "environment.sv"
`include "test.sv"

endpackage
